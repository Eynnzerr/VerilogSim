module reg74HC374(
	input OE,CP,[7:0]D,
	output reg[7:0]Q
);
	
	
endmodule